module mem_main(

);






endmodule