module mux_three_to_one(

);






endmodule