module reg_pipe_stage_a(
	input wire	[15:0] in

);






endmodule