module reg_pipe_stage_b(

);






endmodule