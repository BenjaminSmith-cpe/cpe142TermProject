module reg_program_counter(
	input wire address[15:0]
);





endmodule