module shift_two(

);






endmodule