module comparator(

);






endmodule