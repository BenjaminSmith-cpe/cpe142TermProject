module pc_adder(

);






endmodule