module jump_adder(

);






endmodule