module sign_extender(

);






endmodule