import types_pkg::*;
import alu_pkg::*;

module top (
	input wire clk,
	input wire rst
);
	
stage_one st1(
	);

stage_two st2(
	);

endmodule
