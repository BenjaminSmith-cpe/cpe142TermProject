module mux_two_to_one(

);






endmodule