module mem_program(

);






endmodule