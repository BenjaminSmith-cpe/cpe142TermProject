module control_main(

);






endmodule