module control_alu(

);






endmodule