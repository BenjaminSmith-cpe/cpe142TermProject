module jump_control(

);






endmodule