module reg_pipe_stage_a(

);






endmodule