package reg_program_counter_pkg